** sch_path: /home/scholes33/Projects/PreLayout/Xschem/readsnm.sch
**.subckt readsnm
XM1 VCC qb1 q1 VCC sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad=0.1218 as=0.1218 pd=1.42 ps=1.42 nrd=0.69047619047619
+ nrs=0.69047619047619 sa=0 sb=0 sd=0 mult=1 m=1
XM2 GND qb1 q1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 ad=0.2436 as=0.2436 pd=2.26 ps=2.26 nrd=0.345238095238095
+ nrs=0.345238095238095 sa=0 sb=0 sd=0 mult=1 m=1
XM3 qb2 q2 VCC VCC sky130_fd_pr__pfet_01v8 L=0.15 W=0.42 nf=1 ad=0.1218 as=0.1218 pd=1.42 ps=1.42 nrd=0.69047619047619
+ nrs=0.69047619047619 sa=0 sb=0 sd=0 mult=1 m=1
XM4 qb2 q2 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.84 nf=1 ad=0.2436 as=0.2436 pd=2.26 ps=2.26 nrd=0.345238095238095
+ nrs=0.345238095238095 sa=0 sb=0 sd=0 mult=1 m=1
XM5 q1 VCC VCC GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad=0.1218 as=0.1218 pd=1.42 ps=1.42 nrd=0.69047619047619
+ nrs=0.69047619047619 sa=0 sb=0 sd=0 mult=1 m=1
XM6 VCC VCC qb2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 nf=1 ad=0.1218 as=0.1218 pd=1.42 ps=1.42 nrd=0.69047619047619
+ nrs=0.69047619047619 sa=0 sb=0 sd=0 mult=1 m=1
V2 q2 GND 1.8V
V1 qb1 GND 1.8V
VCC VCC GND {supl}
**** begin user architecture code

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.param temp=27
.param supl=1.8

.dc V1 0 1.8 0.01 V2 0 1.8 0.01
.control
run
setplot
setplot dc1
plot q1 vs qb1 q2 vs qb2
wrdata /home/scholes33/Projects/PreLayout/Xschem/readsnm.txt q1 qb1 q2 qb2
.endc
.end


**** end user architecture code
**.ends
.GLOBAL GND
.end