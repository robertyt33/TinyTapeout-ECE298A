magic
tech sky130A
timestamp 1764124684
<< nwell >>
rect 652 1416 950 1542
<< nmos >>
rect 738 1222 756 1306
rect 870 1222 888 1306
rect 696 1090 738 1114
rect 840 1090 882 1114
<< pmos >>
rect 738 1434 756 1476
rect 870 1434 888 1476
<< ndiff >>
rect 696 1298 738 1306
rect 696 1230 702 1298
rect 720 1230 738 1298
rect 696 1222 738 1230
rect 756 1298 798 1306
rect 756 1230 774 1298
rect 792 1230 798 1298
rect 756 1222 798 1230
rect 828 1298 870 1306
rect 828 1230 834 1298
rect 852 1230 870 1298
rect 828 1222 870 1230
rect 888 1298 930 1306
rect 888 1230 906 1298
rect 924 1230 930 1298
rect 888 1222 930 1230
rect 696 1144 738 1150
rect 696 1126 705 1144
rect 729 1126 738 1144
rect 696 1114 738 1126
rect 840 1144 882 1150
rect 840 1126 849 1144
rect 873 1126 882 1144
rect 840 1114 882 1126
rect 696 1078 738 1090
rect 696 1060 705 1078
rect 729 1060 738 1078
rect 696 1054 738 1060
rect 840 1078 882 1090
rect 840 1060 849 1078
rect 873 1060 882 1078
rect 840 1054 882 1060
<< pdiff >>
rect 696 1468 738 1476
rect 696 1442 702 1468
rect 720 1442 738 1468
rect 696 1434 738 1442
rect 756 1468 798 1476
rect 756 1442 774 1468
rect 792 1442 798 1468
rect 756 1434 798 1442
rect 828 1468 870 1476
rect 828 1442 834 1468
rect 852 1442 870 1468
rect 828 1434 870 1442
rect 888 1468 930 1476
rect 888 1442 906 1468
rect 924 1442 930 1468
rect 888 1434 930 1442
<< ndiffc >>
rect 702 1230 720 1298
rect 774 1230 792 1298
rect 834 1230 852 1298
rect 906 1230 924 1298
rect 705 1126 729 1144
rect 849 1126 873 1144
rect 705 1060 729 1078
rect 849 1060 873 1078
<< pdiffc >>
rect 702 1442 720 1468
rect 774 1442 792 1468
rect 834 1442 852 1468
rect 906 1442 924 1468
<< psubdiff >>
rect 698 1178 738 1195
rect 764 1178 812 1195
rect 834 1178 878 1195
<< nsubdiff >>
rect 700 1523 877 1524
rect 700 1506 726 1523
rect 756 1506 804 1523
rect 834 1506 877 1523
rect 700 1504 877 1506
<< psubdiffcont >>
rect 738 1178 764 1195
rect 812 1178 834 1195
<< nsubdiffcont >>
rect 726 1506 756 1523
rect 804 1506 834 1523
<< poly >>
rect 738 1476 756 1494
rect 870 1476 888 1494
rect 738 1406 756 1434
rect 814 1406 846 1414
rect 738 1388 821 1406
rect 839 1388 846 1406
rect 738 1306 756 1388
rect 814 1380 846 1388
rect 814 1350 846 1358
rect 870 1350 888 1434
rect 814 1332 821 1350
rect 839 1332 888 1350
rect 814 1324 846 1332
rect 870 1306 888 1332
rect 738 1208 756 1222
rect 870 1208 888 1222
rect 770 1114 808 1118
rect 678 1090 696 1114
rect 738 1112 840 1114
rect 738 1094 778 1112
rect 800 1094 840 1112
rect 738 1090 840 1094
rect 882 1090 900 1114
rect 770 1086 808 1090
<< polycont >>
rect 821 1388 839 1406
rect 821 1332 839 1350
rect 778 1094 800 1112
<< locali >>
rect 696 1524 882 1528
rect 696 1507 703 1524
rect 720 1523 882 1524
rect 720 1507 726 1523
rect 696 1506 726 1507
rect 756 1506 804 1523
rect 834 1506 840 1523
rect 857 1506 882 1523
rect 696 1500 882 1506
rect 702 1476 720 1500
rect 834 1476 852 1500
rect 696 1468 726 1476
rect 696 1442 702 1468
rect 720 1442 726 1468
rect 696 1434 726 1442
rect 768 1468 798 1476
rect 768 1442 774 1468
rect 792 1442 798 1468
rect 768 1434 798 1442
rect 828 1468 858 1476
rect 828 1442 834 1468
rect 852 1442 858 1468
rect 828 1434 858 1442
rect 900 1468 930 1476
rect 900 1442 906 1468
rect 924 1442 930 1468
rect 900 1434 930 1442
rect 774 1374 792 1434
rect 814 1406 846 1414
rect 906 1406 924 1434
rect 814 1388 821 1406
rect 839 1388 924 1406
rect 814 1380 846 1388
rect 660 1356 792 1374
rect 660 1144 678 1356
rect 774 1350 792 1356
rect 814 1350 846 1358
rect 774 1332 821 1350
rect 839 1332 846 1350
rect 774 1306 792 1332
rect 814 1324 846 1332
rect 906 1306 924 1388
rect 696 1298 726 1306
rect 696 1230 702 1298
rect 720 1230 726 1298
rect 696 1222 726 1230
rect 768 1298 798 1306
rect 768 1230 774 1298
rect 792 1230 798 1298
rect 768 1222 798 1230
rect 828 1298 858 1306
rect 828 1230 834 1298
rect 852 1230 858 1298
rect 828 1222 858 1230
rect 900 1298 930 1306
rect 900 1230 906 1298
rect 924 1230 930 1298
rect 900 1222 930 1230
rect 702 1198 720 1222
rect 834 1198 852 1222
rect 696 1195 882 1198
rect 696 1178 702 1195
rect 724 1178 738 1195
rect 764 1178 812 1195
rect 834 1178 838 1195
rect 860 1178 882 1195
rect 696 1175 882 1178
rect 696 1144 738 1150
rect 660 1126 705 1144
rect 729 1126 738 1144
rect 696 1120 738 1126
rect 840 1144 882 1150
rect 906 1144 924 1222
rect 840 1126 849 1144
rect 873 1126 924 1144
rect 840 1120 882 1126
rect 770 1112 808 1118
rect 770 1092 776 1112
rect 802 1092 808 1112
rect 770 1086 808 1092
rect 652 1080 674 1084
rect 696 1080 738 1084
rect 652 1062 656 1080
rect 674 1078 738 1080
rect 674 1062 705 1078
rect 652 1056 674 1062
rect 696 1060 705 1062
rect 729 1060 738 1078
rect 696 1054 738 1060
rect 840 1080 882 1084
rect 906 1080 928 1084
rect 840 1078 910 1080
rect 840 1060 849 1078
rect 873 1062 910 1078
rect 873 1060 882 1062
rect 840 1054 882 1060
rect 906 1056 928 1062
<< viali >>
rect 703 1507 720 1524
rect 840 1506 857 1523
rect 702 1178 724 1195
rect 838 1178 860 1195
rect 776 1094 778 1112
rect 778 1094 800 1112
rect 800 1094 802 1112
rect 776 1092 802 1094
rect 656 1062 674 1080
rect 910 1062 928 1080
<< metal1 >>
rect 652 1080 680 1578
rect 696 1524 766 1528
rect 696 1507 703 1524
rect 720 1507 766 1524
rect 696 1500 766 1507
rect 796 1523 882 1528
rect 796 1506 840 1523
rect 857 1506 882 1523
rect 796 1500 882 1506
rect 696 1201 882 1204
rect 696 1195 771 1201
rect 696 1178 702 1195
rect 724 1178 771 1195
rect 696 1175 771 1178
rect 805 1195 882 1201
rect 805 1178 838 1195
rect 860 1178 882 1195
rect 805 1175 882 1178
rect 770 1116 808 1118
rect 770 1086 776 1116
rect 802 1086 808 1116
rect 652 1062 656 1080
rect 674 1062 680 1080
rect 652 1054 680 1062
rect 904 1080 932 1578
rect 904 1062 910 1080
rect 928 1062 932 1080
rect 904 1054 932 1062
<< via1 >>
rect 766 1500 796 1528
rect 771 1175 805 1201
rect 776 1112 802 1116
rect 776 1092 802 1112
rect 776 1086 802 1092
<< metal2 >>
rect 652 1500 766 1528
rect 796 1500 950 1528
rect 652 1201 950 1204
rect 652 1175 771 1201
rect 805 1175 950 1201
rect 652 1174 950 1175
rect 770 1116 808 1118
rect 770 1114 776 1116
rect 652 1090 776 1114
rect 770 1086 776 1090
rect 802 1114 808 1116
rect 802 1090 950 1114
rect 802 1086 808 1090
<< labels >>
rlabel locali 906 1388 924 1406 1 qbar
port 4 n
rlabel locali 660 1356 678 1374 1 q
port 6 n
rlabel locali 666 1062 684 1080 1 bl
port 2 n
rlabel metal2 696 1175 882 1204 1 gnd
port 9 n
rlabel locali 894 1062 912 1080 1 blbar
port 3 n
rlabel nwell 696 1500 882 1528 1 vdd
port 8 n
rlabel metal2 770 1086 808 1118 1 wl
port 10 n
<< end >>
