magic
tech sky130A
timestamp 1764302968
<< nwell >>
rect -54 108 142 192
<< nmos >>
rect -62 -82 -44 -40
rect 2 -82 20 2
rect 66 -82 84 2
rect 132 -82 150 -40
<< pmos >>
rect 2 126 20 168
rect 66 126 84 168
<< ndiff >>
rect -36 -6 2 2
rect -36 -40 -32 -6
rect -96 -50 -62 -40
rect -96 -74 -92 -50
rect -74 -74 -62 -50
rect -96 -82 -62 -74
rect -44 -74 -32 -40
rect -14 -74 2 -6
rect -44 -82 2 -74
rect 20 -6 66 2
rect 20 -74 32 -6
rect 50 -74 66 -6
rect 20 -82 66 -74
rect 84 -6 124 2
rect 84 -74 98 -6
rect 116 -40 124 -6
rect 116 -74 132 -40
rect 84 -82 132 -74
rect 150 -48 184 -40
rect 150 -74 162 -48
rect 180 -74 184 -48
rect 150 -82 184 -74
<< pdiff >>
rect -36 160 2 168
rect -36 134 -32 160
rect -14 134 2 160
rect -36 126 2 134
rect 20 160 66 168
rect 20 134 32 160
rect 50 134 66 160
rect 20 126 66 134
rect 84 160 124 168
rect 84 134 98 160
rect 116 134 124 160
rect 84 126 124 134
<< ndiffc >>
rect -92 -74 -74 -50
rect -32 -74 -14 -6
rect 32 -74 50 -6
rect 98 -74 116 -6
rect 162 -74 180 -48
<< pdiffc >>
rect -32 134 -14 160
rect 32 134 50 160
rect 98 134 116 160
<< poly >>
rect 2 168 20 186
rect 66 168 84 186
rect 2 102 20 126
rect 2 96 44 102
rect 2 78 18 96
rect 36 78 44 96
rect 2 72 44 78
rect 2 2 20 72
rect 66 50 84 126
rect 42 44 84 50
rect 42 26 50 44
rect 68 26 84 44
rect 42 20 84 26
rect 66 2 84 20
rect -62 -40 -44 -26
rect 132 -40 150 -26
rect -62 -128 -44 -82
rect 2 -96 20 -82
rect 66 -96 84 -82
rect 132 -128 150 -82
rect -62 -138 -22 -128
rect -62 -156 -48 -138
rect -30 -156 -22 -138
rect -62 -164 -22 -156
rect 110 -138 150 -128
rect 110 -156 118 -138
rect 136 -156 150 -138
rect 110 -164 150 -156
rect -62 -166 -42 -164
rect 132 -166 150 -164
<< polycont >>
rect 18 78 36 96
rect 50 26 68 44
rect -48 -156 -30 -138
rect 118 -156 136 -138
<< locali >>
rect 28 176 34 194
rect 52 176 58 194
rect -36 160 -6 168
rect -36 134 -32 160
rect -14 134 -6 160
rect -36 126 -6 134
rect 28 160 58 176
rect 28 134 32 160
rect 50 134 58 160
rect 28 126 58 134
rect 94 160 124 168
rect 94 134 98 160
rect 116 134 124 160
rect 94 126 124 134
rect -30 38 -12 126
rect 100 102 118 126
rect 10 96 118 102
rect 10 78 18 96
rect 36 84 118 96
rect 36 78 44 84
rect 10 72 44 78
rect 42 44 76 50
rect 42 38 50 44
rect -30 26 50 38
rect 68 26 76 44
rect -30 20 76 26
rect -30 2 -12 20
rect 100 2 118 84
rect -36 -6 -6 2
rect -96 -48 -70 -40
rect -96 -74 -92 -48
rect -74 -74 -70 -48
rect -96 -82 -70 -74
rect -36 -74 -32 -6
rect -14 -74 -6 -6
rect -36 -82 -6 -74
rect 28 -6 58 2
rect 28 -74 32 -6
rect 50 -74 58 -6
rect 28 -92 58 -74
rect 94 -6 124 2
rect 94 -74 98 -6
rect 116 -74 124 -6
rect 94 -82 124 -74
rect 158 -48 184 -40
rect 158 -74 162 -48
rect 180 -74 184 -48
rect 158 -82 184 -74
rect 28 -110 32 -92
rect 54 -110 58 -92
rect 28 -114 58 -110
rect -56 -138 -22 -128
rect -56 -156 -48 -138
rect -30 -156 -22 -138
rect -56 -164 -22 -156
rect 110 -138 144 -128
rect 110 -156 118 -138
rect 136 -156 144 -138
rect 110 -164 144 -156
<< viali >>
rect 34 176 52 194
rect -92 -50 -74 -48
rect -92 -74 -74 -50
rect 162 -74 180 -48
rect 32 -110 54 -92
rect -48 -156 -30 -138
rect 118 -156 136 -138
<< metal1 >>
rect -96 -48 -70 212
rect 24 172 30 198
rect 56 172 62 198
rect -96 -74 -92 -48
rect -74 -74 -70 -48
rect -96 -166 -70 -74
rect 158 -48 184 212
rect 158 -74 162 -48
rect 180 -74 184 -48
rect 26 -84 60 -82
rect 26 -110 30 -84
rect 56 -110 60 -84
rect 26 -114 60 -110
rect -56 -132 -20 -128
rect -56 -162 -48 -132
rect -22 -162 -20 -132
rect -56 -166 -20 -162
rect 108 -132 144 -128
rect 108 -162 110 -132
rect 136 -162 144 -132
rect 108 -166 144 -162
rect 158 -166 184 -74
<< via1 >>
rect 30 194 56 198
rect 30 176 34 194
rect 34 176 52 194
rect 52 176 56 194
rect 30 172 56 176
rect 30 -92 56 -84
rect 30 -110 32 -92
rect 32 -110 54 -92
rect 54 -110 56 -92
rect -48 -138 -22 -132
rect -48 -156 -30 -138
rect -30 -156 -22 -138
rect -48 -162 -22 -156
rect 110 -138 136 -132
rect 110 -156 118 -138
rect 118 -156 136 -138
rect 110 -162 136 -156
<< metal2 >>
rect -96 172 30 198
rect 56 172 184 198
rect 26 -84 100 -82
rect 26 -110 30 -84
rect 56 -110 62 -84
rect 26 -112 62 -110
rect 90 -112 100 -84
rect 26 -114 100 -112
rect -96 -132 184 -128
rect -96 -162 -48 -132
rect -22 -162 110 -132
rect 136 -162 184 -132
rect -96 -166 184 -162
<< via2 >>
rect 62 -112 90 -84
<< metal3 >>
rect 26 -82 114 -80
rect -96 -84 184 -82
rect -96 -112 62 -84
rect 90 -112 184 -84
rect -96 -116 184 -112
<< labels >>
rlabel locali 10 72 44 102 1 qbar
port 1 n
rlabel metal1 -96 -82 -70 -40 1 bl
port 3 n
rlabel metal1 158 -82 184 -40 1 blbar
port 4 n
rlabel locali 42 20 76 50 1 q
port 2 n
rlabel metal2 16 -164 70 -128 1 wl
port 5 n
rlabel metal2 26 174 62 198 1 vdd
port 6 n
rlabel metal3 26 -112 60 -82 1 gnd
port 7 n
<< end >>
