* NGSPICE file created from 6T_SRAM_1bit_Type1b.ext - technology: sky130A

.subckt x6T_SRAM_1bit_Type1b qbar q bl blbar wl vdd gnd
X0 blbar wl qbar SUB sky130_fd_pr__nfet_01v8 ad=0.1428 pd=1.52 as=0.1848 ps=1.32 w=0.42 l=0.18
X1 q wl bl SUB sky130_fd_pr__nfet_01v8 ad=0.1764 pd=1.3 as=0.1428 ps=1.52 w=0.42 l=0.18
X2 qbar q gnd SUB sky130_fd_pr__nfet_01v8 ad=0.1848 pd=1.32 as=0.1932 ps=1.3 w=0.84 l=0.18
X3 gnd qbar q SUB sky130_fd_pr__nfet_01v8 ad=0.1932 pd=1.3 as=0.1764 ps=1.3 w=0.84 l=0.18
X4 qbar q vdd w_n54_108# sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.64 as=0.0966 ps=0.88 w=0.42 l=0.18
X5 vdd qbar q w_n54_108# sky130_fd_pr__pfet_01v8 ad=0.0966 pd=0.88 as=0.1596 ps=1.6 w=0.42 l=0.18
C0 qbar blbar 0.06872f
C1 bl w_n54_108# 0.00579f
C2 wl q 0.03298f
C3 q gnd 0.11079f
C4 wl gnd 0.20082f
C5 vdd bl 0.05123f
C6 q blbar 0.0161f
C7 qbar bl 0.01658f
C8 wl blbar 0.09277f
C9 blbar gnd 0.03697f
C10 vdd w_n54_108# 0.02115f
C11 qbar w_n54_108# 0.04742f
C12 q bl 0.06839f
C13 wl bl 0.09277f
C14 qbar vdd 0.07319f
C15 bl gnd 0.03519f
C16 bl blbar 0.04942f
C17 q w_n54_108# 0.03965f
C18 wl w_n54_108# 0.00595f
C19 w_n54_108# gnd 0.00317f
C20 w_n54_108# blbar 0.00585f
C21 q vdd 0.0486f
C22 wl vdd 0.03392f
C23 qbar q 0.25781f
C24 qbar wl 0.03393f
C25 vdd gnd 0.0268f
C26 qbar gnd 0.07836f
C27 vdd blbar 0.05105f
C28 blbar SUB 0.26304f
C29 gnd SUB 0.30417f
C30 bl SUB 0.26292f
C31 wl SUB 0.67354f
C32 vdd SUB 0.19783f
C33 q SUB 0.35241f
C34 qbar SUB 0.34852f
C35 w_n54_108# SUB 0.19757f
.ends

